library verilog;
use verilog.vl_types.all;
entity sistema_vlg_vec_tst is
end sistema_vlg_vec_tst;
